module half_sub
