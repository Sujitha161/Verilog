module tb_dcon;
	reg d,clk,rst;
	wire q;
cd uut (.d(d),.clk(clk),.rst(rst),.q(q));
	always #5 clk = ~clk;
	initial begin 
		clk=1;rst=0;d=0;
		#10;
		d=1;
		#10;rst=1;d=0;#10;
		d=1;#5 ;rst=0;#10;d=1;
		#100 $finish;
	end
	initial begin
	       $dumpfile("out_dcon.vcd");
       	       $dumpvars(0,tb_dcon);
	       $monitor("time=%0t,d=%b,clk=%b,rst=%b,q=%b",$time,d,clk,rst,q);
       end
       endmodule

